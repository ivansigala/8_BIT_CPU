
//Diego Iván Sigala Sánchez
//Sistemas digitales

module ROM(
    input [7:0]addr,
    output reg [11:0]out
    );
    
    
    always @ (*) begin
        case(addr)
            1: out = 12'hF00;
            2: out = 12'h500;
            3: out = 12'hF00;
            4: out = 12'h501;
            5: out = 12'hF05;
            6: out = 12'h201;
            7: out = 12'h001;
            8: out = 12'h101;
            9: out = 12'h501;
            10: out = 12'h000;
            11: out = 12'h700;
            12: out = 12'h605;
            13: out = 12'h001;
            14: out = 12'h9FF;
            15: out = 12'h9FF;
            16: out = 12'h9FF;
            17: out = 12'h9FF;
            18: out = 12'h9FF;
            19: out = 12'h9FF;
            20: out = 12'h9FF;
            21: out = 12'h9FF;
            22: out = 12'h9FF;
            23: out = 12'h9FF;
            24: out = 12'h9FF;
            25: out = 12'h9FF;
            26: out = 12'h9FF;
            27: out = 12'h9FF;
            28: out = 12'h9FF;
            29: out = 12'h9FF;
            30: out = 12'h9FF;
            31: out = 12'h9FF;
            32: out = 12'h9FF;
            33: out = 12'h9FF;
            34: out = 12'h9FF;
            35: out = 12'h9FF;
            36: out = 12'h9FF;
            37: out = 12'h9FF;
            38: out = 12'h9FF;
            39: out = 12'h9FF;
            40: out = 12'h9FF;
            41: out = 12'h9FF;
            42: out = 12'h9FF;
            43: out = 12'h9FF;
            44: out = 12'h9FF;
            45: out = 12'h9FF;
            46: out = 12'h9FF;
            47: out = 12'h9FF;
            48: out = 12'h9FF;
            49: out = 12'h9FF;
            50: out = 12'h9FF;
            51: out = 12'h9FF;
            52: out = 12'h9FF;
            53: out = 12'h9FF;
            54: out = 12'h9FF;
            55: out = 12'h9FF;
            56: out = 12'h9FF;
            57: out = 12'h9FF;
            58: out = 12'h9FF;
            59: out = 12'h9FF;
            60: out = 12'h9FF;
            61: out = 12'h9FF;
            62: out = 12'h9FF;
            63: out = 12'h9FF;
            64: out = 12'h9FF;
            65: out = 12'h9FF;
            66: out = 12'h9FF;
            67: out = 12'h9FF;
            68: out = 12'h9FF;
            69: out = 12'h9FF;
            70: out = 12'h9FF;
            71: out = 12'h9FF;
            72: out = 12'h9FF;
            73: out = 12'h9FF;
            74: out = 12'h9FF;
            75: out = 12'h9FF;
            76: out = 12'h9FF;
            77: out = 12'h9FF;
            78: out = 12'h9FF;
            79: out = 12'h9FF;
            80: out = 12'h9FF;
            81: out = 12'h9FF;
            82: out = 12'h9FF;
            83: out = 12'h9FF;
            84: out = 12'h9FF;
            85: out = 12'h9FF;
            86: out = 12'h9FF;
            87: out = 12'h9FF;
            88: out = 12'h9FF;
            89: out = 12'h9FF;
            90: out = 12'h9FF;
            91: out = 12'h9FF;
            92: out = 12'h9FF;
            93: out = 12'h9FF;
            94: out = 12'h9FF;
            95: out = 12'h9FF;
            96: out = 12'h9FF;
            97: out = 12'h9FF;
            98: out = 12'h9FF;
            99: out = 12'h9FF;
            100: out = 12'h9FF;
            101: out = 12'h9FF;
            102: out = 12'h9FF;
            103: out = 12'h9FF;
            104: out = 12'h9FF;
            105: out = 12'h9FF;
            106: out = 12'h9FF;
            107: out = 12'h9FF;
            108: out = 12'h9FF;
            109: out = 12'h9FF;
            110: out = 12'h9FF;
            111: out = 12'h9FF;
            112: out = 12'h9FF;
            113: out = 12'h9FF;
            114: out = 12'h9FF;
            115: out = 12'h9FF;
            116: out = 12'h9FF;
            117: out = 12'h9FF;
            118: out = 12'h9FF;
            119: out = 12'h9FF;
            120: out = 12'h9FF;
            121: out = 12'h9FF;
            122: out = 12'h9FF;
            123: out = 12'h9FF;
            124: out = 12'h9FF;
            125: out = 12'h9FF;
            126: out = 12'h9FF;
            127: out = 12'h9FF;
            128: out = 12'h9FF;
            129: out = 12'h9FF;
            130: out = 12'h9FF;
            131: out = 12'h9FF;
            132: out = 12'h9FF;
            133: out = 12'h9FF;
            134: out = 12'h9FF;
            135: out = 12'h9FF;
            136: out = 12'h9FF;
            137: out = 12'h9FF;
            138: out = 12'h9FF;
            139: out = 12'h9FF;
            140: out = 12'h9FF;
            141: out = 12'h9FF;
            142: out = 12'h9FF;
            143: out = 12'h9FF;
            144: out = 12'h9FF;
            145: out = 12'h9FF;
            146: out = 12'h9FF;
            147: out = 12'h9FF;
            148: out = 12'h9FF;
            149: out = 12'h9FF;
            150: out = 12'h9FF;
            151: out = 12'h9FF;
            152: out = 12'h9FF;
            153: out = 12'h9FF;
            154: out = 12'h9FF;
            155: out = 12'h9FF;
            156: out = 12'h9FF;
            157: out = 12'h9FF;
            158: out = 12'h9FF;
            159: out = 12'h9FF;
            160: out = 12'h9FF;
            161: out = 12'h9FF;
            162: out = 12'h9FF;
            163: out = 12'h9FF;
            164: out = 12'h9FF;
            165: out = 12'h9FF;
            166: out = 12'h9FF;
            167: out = 12'h9FF;
            168: out = 12'h9FF;
            169: out = 12'h9FF;
            170: out = 12'h9FF;
            171: out = 12'h9FF;
            172: out = 12'h9FF;
            173: out = 12'h9FF;
            174: out = 12'h9FF;
            175: out = 12'h9FF;
            176: out = 12'h9FF;
            177: out = 12'h9FF;
            178: out = 12'h9FF;
            179: out = 12'h9FF;
            180: out = 12'h9FF;
            181: out = 12'h9FF;
            182: out = 12'h9FF;
            183: out = 12'h9FF;
            184: out = 12'h9FF;
            185: out = 12'h9FF;
            186: out = 12'h9FF;
            187: out = 12'h9FF;
            188: out = 12'h9FF;
            189: out = 12'h9FF;
            190: out = 12'h9FF;
            191: out = 12'h9FF;
            192: out = 12'h9FF;
            193: out = 12'h9FF;
            194: out = 12'h9FF;
            195: out = 12'h9FF;
            196: out = 12'h9FF;
            197: out = 12'h9FF;
            198: out = 12'h9FF;
            199: out = 12'h9FF;
            200: out = 12'h9FF;
            201: out = 12'h9FF;
            202: out = 12'h9FF;
            203: out = 12'h9FF;
            204: out = 12'h9FF;
            205: out = 12'h9FF;
            206: out = 12'h9FF;
            207: out = 12'h9FF;
            208: out = 12'h9FF;
            209: out = 12'h9FF;
            210: out = 12'h9FF;
            211: out = 12'h9FF;
            212: out = 12'h9FF;
            213: out = 12'h9FF;
            214: out = 12'h9FF;
            215: out = 12'h9FF;
            216: out = 12'h9FF;
            217: out = 12'h9FF;
            218: out = 12'h9FF;
            219: out = 12'h9FF;
            220: out = 12'h9FF;
            221: out = 12'h9FF;
            222: out = 12'h9FF;
            223: out = 12'h9FF;
            224: out = 12'h9FF;
            225: out = 12'h9FF;
            226: out = 12'h9FF;
            227: out = 12'h9FF;
            228: out = 12'h9FF;
            229: out = 12'h9FF;
            230: out = 12'h9FF;
            231: out = 12'h9FF;
            232: out = 12'h9FF;
            233: out = 12'h9FF;
            234: out = 12'h9FF;
            235: out = 12'h9FF;
            236: out = 12'h9FF;
            237: out = 12'h9FF;
            238: out = 12'h9FF;
            239: out = 12'h9FF;
            240: out = 12'h9FF;
            241: out = 12'h9FF;
            242: out = 12'h9FF;
            243: out = 12'h9FF;
            244: out = 12'h9FF;
            245: out = 12'h9FF;
            246: out = 12'h9FF;
            247: out = 12'h9FF;
            248: out = 12'h9FF;
            249: out = 12'h9FF;
            250: out = 12'h9FF;
            251: out = 12'h9FF;
            252: out = 12'h9FF;
            253: out = 12'h9FF;
            254: out = 12'h9FF;
            255: out = 12'h9FF;
        endcase
    end

    
endmodule
